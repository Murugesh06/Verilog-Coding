`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.08.2025 15:24:56
// Design Name: 
// Module Name: function_sum_of_2numbers
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module function_sum_of_2numbers;
function [7:0]sum;
input [7:0]a,b;
begin
sum=a+b;
end
endfunction
endmodule
